core_tlib